LIBRARY ieee;
USE ieee.std_logic_1164.all;
library digital_components;
use digital_components.fullAdder_v1_package.all;

ENTITY RippleCarryAdder IS 
  PORT (A, B          : IN  STD_LOGIC_vector(3 downto 0);
        s             : out std_logic_vector(3 downto 0);
        c             : out STD_LOGIC);
END RippleCarryAdder;

architecture structural of RippleCarryAdder is
signal ripple_carry : std_logic_vector(3 downto 0); 
--signal c1, c2, c3;
begin 

--fullAdder0  : fullAdder port map (A(0),  B(0),  '0',             ripple_carry(0), s(0));
--fullAdder1  : fullAdder port map (A(1),  B(1),  ripple_carry(0), ripple_carry(1), s(1));
--fullAdder2  : fullAdder port map (A(2),  B(2),  ripple_carry(1), ripple_carry(2), s(2));
--fullAdder3  : fullAdder port map (A(3),  B(3),  ripple_carry(2), c,               s(3));

fullAdder1  : fullAdder_v1_structure port map (A(0),  B(0),  '0',               ripple_carry(0), s(0));
  G1: for i in 1 to 3 generate
         fullAdders  : fullAdder_v1_structure port map (A(i),  B(i),  ripple_carry(i-1), ripple_carry(i), s(i));
  end generate;
c <= ripple_carry(3);

end structural;
