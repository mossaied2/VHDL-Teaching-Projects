-- Testbench for OR gate
library IEEE;
use IEEE.std_logic_1164.all;
USE ieee.std_logic_unsigned.all ;

entity comparatorNbits_v3_structure_testbench is
-- empty
end comparatorNbits_v3_structure_testbench; 

architecture comparatorNbits_v3_structure_tb of comparatorNbits_v3_structure_testbench is

-- DUT component
component comparatorNbits_v3_structure is
PORT (A, B  : IN STD_LOGIC_vector(15 downto 0);
AeqB, AltB, AgtB  : OUT STD_LOGIC);
end component;

signal AeqB_out, AltB_out, AgtB_out : std_logic;
signal A_in, B_in : std_logic_vector(15 downto 0);

begin

  -- Connect DUT
  DUT: comparatorNbits_v3_structure port map(A_in, B_in, AeqB_out, AltB_out, AgtB_out);

  process
  begin

    A_in <= x"0011";
    B_in <= x"0001";
    wait for 1 ns;
     
    A_in <= x"0010";
    B_in <= x"0101";
    wait for 1 ns;
     
    A_in <= x"f111";
    B_in <= x"1f11";
    wait for 1 ns;
     
    A_in <= x"0110";
    B_in <= x"1000";
    wait for 1 ns;
    
    A_in <= x"0000";
    B_in <= x"0000";
    wait for 1 ns;
  

A_in <= x"0011";
    B_in <= x"0001";
    wait for 1 ns;
     
    A_in <= x"0010";
    B_in <= x"0101";
    wait for 1 ns;
     
    A_in <= x"f111";
    B_in <= x"1f11";
    wait for 1 ns;
     
    A_in <= x"0110";
    B_in <= x"1000";
    wait for 1 ns;
    
    A_in <= x"0000";
    B_in <= x"0000";
    wait for 1 ns;
    assert false report "Test done." severity note;
    wait;
  end process;
end comparatorNbits_v3_structure_tb;

