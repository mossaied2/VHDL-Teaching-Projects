-- Testbench for OR gate
library IEEE;
use IEEE.std_logic_1164.all;
 
entity JK_FF_testbench is
-- empty
end JK_FF_testbench; 

architecture JK_FF_tb of JK_FF_testbench is

-- DUT component
component JK_FF is
  PORT (j, k, clk, reset   : IN  STD_LOGIC;
        Q, Q_bar           : out  STD_LOGIC);
end component;

signal j_in, k_in : STD_LOGIC;
signal clk_in : std_logic := '0';
signal reset_in : std_logic := '1';
signal Q_out : STD_LOGIC ;
signal Q_bar_out : STD_LOGIC ;

begin

  -- Connect DUT
  DUT: JK_FF port map(j_in, k_in, clk_in, reset_in, Q_out, Q_bar_out);

  -- Process for generating the clock
  clk_in <= not clk_in after 1.010 ns;

  process
  begin
    j_in <= '1';reset_in <= '1';
    k_in <= '0';
    wait for 1 ns; 
    j_in <= '1';reset_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';reset_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;  
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;  
  j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;   
 j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;   
 j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;  
  j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;  
  j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;    
j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;    
j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;   
 j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '1';
    wait for 1 ns; 
    j_in <= '0';
    k_in <= '1';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '0';
    k_in <= '0';
    wait for 1 ns;
    j_in <= '1';
    k_in <= '0';
    wait for 1 ns;
    
    assert false report "Test done." severity note;
    wait;
  end process;
end JK_FF_tb;

